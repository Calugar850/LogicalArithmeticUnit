----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 21.11.2021 14:48:46
-- Design Name: 
-- Module Name: unitate_conversie_in_C2 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity unitate_conversie_in_C2 is
  Port (Yin : in std_logic_vector (7 downto 0);
        Yout : out std_logic_vector (7 downto 0));
end unitate_conversie_in_C2;

architecture Behavioral of unitate_conversie_in_C2 is

begin

Yout<=(not Yin) + '1';
end Behavioral;
